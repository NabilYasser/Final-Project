module Serializer_Top (
    input wire Ser_En,
    input wire RST,
    input wire clk,
    input wire Data_Valid,
    input wire [7:0] P_Data_Top,
    output wire Ser_Data_Top,
    output wire Ser_Done

);
wire [2:0] Counter_Top;
//wire Counter_RST= Ser_En & RST;

Counter u_Counter(
    .RST     (RST     ),
    .clk     (clk     ),
    .Counter (Counter_Top ),
    .Ser_En  (Ser_En) ,
    .Finish  (Ser_Done  )
);

Serializer u_Serializer(
    .P_Data   (P_Data_Top   ),
    .clk      (clk      ),
    .rst(RST),
    .Ser_En(Ser_En),
    .Data_Valid(Data_Valid),
    .Counter  (Counter_Top  ),
    .Ser_Data (Ser_Data_Top )
);


    
endmodule